/*

Copyright (c) 2015 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * AXI4-Stream frame length adjuster
 */
module axis_frame_length_adjust #
(
    parameter DATA_WIDTH = 1,
    parameter KEEP_WIDTH = (DATA_WIDTH/8)
)
(
    input  wire                   clk,
    input  wire                   rst,

    /*
     * AXI input
     */
    input  wire [DATA_WIDTH-1:0]  input_axis_tdata,
    input  wire [KEEP_WIDTH-1:0]  input_axis_tkeep,
    input  wire                   input_axis_tvalid,
    output wire                   input_axis_tready,
    input  wire                   input_axis_tlast,
    input  wire                   input_axis_tuser,

    /*
     * AXI output
     */
    output wire [DATA_WIDTH-1:0]  output_axis_tdata,
    output wire [KEEP_WIDTH-1:0]  output_axis_tkeep,
    output wire                   output_axis_tvalid,
    input  wire                   output_axis_tready,
    output wire                   output_axis_tlast,
    output wire                   output_axis_tuser,

    /*
     * Status
     */
    output wire                   status_valid,
    input  wire                   status_ready,
    output wire                   status_frame_pad,
    output wire                   status_frame_truncate,
    output wire [15:0]            status_frame_length,
    output wire [15:0]            status_frame_original_length,

    /*
     * Configuration
     */
    input  wire [15:0]            length_min,
    input  wire [15:0]            length_max
);

// bus word width
localparam DATA_WORD_WIDTH = DATA_WIDTH / KEEP_WIDTH;

// bus width assertions
initial begin
    if (DATA_WORD_WIDTH * KEEP_WIDTH != DATA_WIDTH) begin
        $error("Error: data width not evenly divisble");
        $finish;
    end
end

// state register
localparam [2:0]
    STATE_IDLE = 3'd0,
    STATE_TRANSFER = 3'd1,
    STATE_PAD = 3'd2,
    STATE_TRUNCATE = 3'd3;

reg [2:0] state_reg = STATE_IDLE, state_next;

// datapath control signals
reg store_last_word;

reg [15:0] frame_ptr_reg = 0, frame_ptr_next;

reg [DATA_WIDTH-1:0] last_word_data_reg = 0;
reg [KEEP_WIDTH-1:0] last_word_keep_reg = 0;

reg last_cycle_tuser_reg = 0, last_cycle_tuser_next;

reg status_valid_reg = 0, status_valid_next;
reg status_frame_pad_reg = 0, status_frame_pad_next;
reg status_frame_truncate_reg = 0, status_frame_truncate_next;
reg [15:0] status_frame_length_reg = 0, status_frame_length_next;
reg [15:0] status_frame_original_length_reg = 0, status_frame_original_length_next;

// internal datapath
reg [DATA_WIDTH-1:0] output_axis_tdata_int;
reg [KEEP_WIDTH-1:0] output_axis_tkeep_int;
reg                  output_axis_tvalid_int;
reg                  output_axis_tready_int = 0;
reg                  output_axis_tlast_int;
reg                  output_axis_tuser_int;
wire                 output_axis_tready_int_early;

reg input_axis_tready_reg = 0, input_axis_tready_next;
assign input_axis_tready = input_axis_tready_reg;

assign status_valid = status_valid_reg;
assign status_frame_pad = status_frame_pad_reg;
assign status_frame_truncate = status_frame_truncate_reg;
assign status_frame_length = status_frame_length_reg;
assign status_frame_original_length = status_frame_original_length_reg;

integer i, word_cnt;

always @* begin
    state_next = STATE_IDLE;

    store_last_word = 0;

    frame_ptr_next = frame_ptr_reg;

    output_axis_tdata_int = 0;
    output_axis_tkeep_int = 0;
    output_axis_tvalid_int = 0;
    output_axis_tlast_int = 0;
    output_axis_tuser_int = 0;

    input_axis_tready_next = 0;

    last_cycle_tuser_next = last_cycle_tuser_reg;

    status_valid_next = status_valid_reg & ~status_ready;
    status_frame_pad_next = status_frame_pad_reg;
    status_frame_truncate_next = status_frame_truncate_reg;
    status_frame_length_next = status_frame_length_reg;
    status_frame_original_length_next = status_frame_original_length_reg;

    case (state_reg)
        STATE_IDLE: begin
            // idle state
            // accept data next cycle if output register ready next cycle
            input_axis_tready_next = output_axis_tready_int_early & (~status_valid_reg | status_ready);

            output_axis_tdata_int = input_axis_tdata;
            output_axis_tkeep_int = input_axis_tkeep;
            output_axis_tvalid_int = input_axis_tvalid;
            output_axis_tlast_int = input_axis_tlast;
            output_axis_tuser_int = input_axis_tuser;

            if (input_axis_tready & input_axis_tvalid) begin
                // transfer through
                word_cnt = 0;
                for (i = 0; i <= KEEP_WIDTH; i = i + 1) begin
                    //bit_cnt = bit_cnt + monitor_axis_tkeep[i];
                    if (input_axis_tkeep == ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-i)) word_cnt = i;
                end
                frame_ptr_next = frame_ptr_reg+word_cnt;

                if (frame_ptr_next >= length_max) begin
                    output_axis_tkeep_int = ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-(length_max - frame_ptr_reg));
                    if (input_axis_tlast) begin
                        status_valid_next = 1;
                        status_frame_pad_next = 0;
                        status_frame_truncate_next = frame_ptr_next > length_max;
                        status_frame_length_next = length_max;
                        status_frame_original_length_next = frame_ptr_next;
                        input_axis_tready_next = output_axis_tready_int_early & status_ready;
                        frame_ptr_next = 0;
                        state_next = STATE_IDLE;
                    end else begin
                        output_axis_tvalid_int = 0;
                        store_last_word = 1;
                        state_next = STATE_TRUNCATE;
                    end
                end else begin
                    if (input_axis_tlast) begin
                        status_frame_original_length_next = frame_ptr_next;
                        if (frame_ptr_next < length_min) begin
                            if (frame_ptr_reg + KEEP_WIDTH < length_min) begin
                                frame_ptr_next = frame_ptr_reg + KEEP_WIDTH;
                                input_axis_tready_next = 0;
                                output_axis_tkeep_int = {KEEP_WIDTH{1'b1}};
                                output_axis_tlast_int = 0;
                                output_axis_tuser_int = 0;
                                last_cycle_tuser_next = input_axis_tuser;
                                state_next = STATE_PAD;
                            end else begin
                                status_valid_next = 1;
                                status_frame_pad_next = 1;
                                status_frame_truncate_next = 0;
                                status_frame_length_next = length_min;
                                input_axis_tready_next = output_axis_tready_int_early & status_ready;
                                output_axis_tkeep_int = ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-(length_min - frame_ptr_reg));
                                frame_ptr_next = 0;
                                state_next = STATE_IDLE;
                            end
                        end else begin
                            status_valid_next = 1;
                            status_frame_pad_next = 0;
                            status_frame_truncate_next = 0;
                            status_frame_length_next = frame_ptr_next;
                            status_frame_original_length_next = frame_ptr_next;
                            input_axis_tready_next = output_axis_tready_int_early & status_ready;
                            frame_ptr_next = 0;
                            state_next = STATE_IDLE;
                        end
                    end else begin
                        state_next = STATE_TRANSFER;
                    end
                end
            end else begin
                state_next = STATE_IDLE;
            end
        end
        STATE_TRANSFER: begin
            // transfer data
            // accept data next cycle if output register ready next cycle
            input_axis_tready_next = output_axis_tready_int_early;

            output_axis_tdata_int = input_axis_tdata;
            output_axis_tkeep_int = input_axis_tkeep;
            output_axis_tvalid_int = input_axis_tvalid;
            output_axis_tlast_int = input_axis_tlast;
            output_axis_tuser_int = input_axis_tuser;

            if (input_axis_tready & input_axis_tvalid) begin
                // transfer through
                word_cnt = 0;
                for (i = 0; i <= KEEP_WIDTH; i = i + 1) begin
                    //bit_cnt = bit_cnt + monitor_axis_tkeep[i];
                    if (input_axis_tkeep == ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-i)) word_cnt = i;
                end
                frame_ptr_next = frame_ptr_reg+word_cnt;

                if (frame_ptr_next >= length_max) begin
                    output_axis_tkeep_int = ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-(length_max - frame_ptr_reg));
                    if (input_axis_tlast) begin
                        status_valid_next = 1;
                        status_frame_pad_next = 0;
                        status_frame_truncate_next = frame_ptr_next > length_max;
                        status_frame_length_next = length_max;
                        status_frame_original_length_next = frame_ptr_next;
                        input_axis_tready_next = output_axis_tready_int_early & status_ready;
                        frame_ptr_next = 0;
                        state_next = STATE_IDLE;
                    end else begin
                        output_axis_tvalid_int = 0;
                        store_last_word = 1;
                        state_next = STATE_TRUNCATE;
                    end
                end else begin
                    if (input_axis_tlast) begin
                        status_frame_original_length_next = frame_ptr_next;
                        if (frame_ptr_next < length_min) begin
                            if (frame_ptr_reg + KEEP_WIDTH < length_min) begin
                                frame_ptr_next = frame_ptr_reg + KEEP_WIDTH;
                                input_axis_tready_next = 0;
                                output_axis_tkeep_int = {KEEP_WIDTH{1'b1}};
                                output_axis_tlast_int = 0;
                                output_axis_tuser_int = 0;
                                last_cycle_tuser_next = input_axis_tuser;
                                state_next = STATE_PAD;
                            end else begin
                                status_valid_next = 1;
                                status_frame_pad_next = 1;
                                status_frame_truncate_next = 0;
                                status_frame_length_next = length_min;
                                input_axis_tready_next = output_axis_tready_int_early & status_ready;
                                output_axis_tkeep_int = ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-(length_min - frame_ptr_reg));
                                frame_ptr_next = 0;
                                state_next = STATE_IDLE;
                            end
                        end else begin
                            status_valid_next = 1;
                            status_frame_pad_next = 0;
                            status_frame_truncate_next = 0;
                            status_frame_length_next = frame_ptr_next;
                            status_frame_original_length_next = frame_ptr_next;
                            input_axis_tready_next = output_axis_tready_int_early & status_ready;
                            frame_ptr_next = 0;
                            state_next = STATE_IDLE;
                        end
                    end else begin
                        state_next = STATE_TRANSFER;
                    end
                end
            end else begin
                state_next = STATE_TRANSFER;
            end
        end
        STATE_PAD: begin
            // pad to minimum length
            input_axis_tready_next = 0;

            output_axis_tdata_int = 0;
            output_axis_tkeep_int = {KEEP_WIDTH{1'b1}};
            output_axis_tvalid_int = 1;
            output_axis_tlast_int = 0;
            output_axis_tuser_int = 0;

            if (output_axis_tready_int) begin
                frame_ptr_next = frame_ptr_reg + KEEP_WIDTH;

                if (frame_ptr_next >= length_min) begin
                    status_valid_next = 1;
                    status_frame_pad_next = 1;
                    status_frame_truncate_next = 0;
                    status_frame_length_next = length_min;
                    input_axis_tready_next = output_axis_tready_int_early & status_ready;
                    output_axis_tkeep_int = ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-(length_min - frame_ptr_reg));
                    output_axis_tlast_int = 1;
                    output_axis_tuser_int = last_cycle_tuser_reg;
                    frame_ptr_next = 0;
                    state_next = STATE_IDLE;
                end else begin
                    state_next = STATE_PAD;
                end
            end else begin
                state_next = STATE_PAD;
            end
        end
        STATE_TRUNCATE: begin
            // drop after maximum length
            input_axis_tready_next = output_axis_tready_int_early;

            output_axis_tdata_int = last_word_data_reg;
            output_axis_tkeep_int = last_word_keep_reg;
            output_axis_tvalid_int = input_axis_tvalid & input_axis_tlast;
            output_axis_tlast_int = input_axis_tlast;
            output_axis_tuser_int = input_axis_tuser;

            if (input_axis_tready & input_axis_tvalid) begin
                word_cnt = 0;
                for (i = 0; i <= KEEP_WIDTH; i = i + 1) begin
                    //bit_cnt = bit_cnt + monitor_axis_tkeep[i];
                    if (input_axis_tkeep == ({KEEP_WIDTH{1'b1}}) >> (KEEP_WIDTH-i)) word_cnt = i;
                end
                frame_ptr_next = frame_ptr_reg+word_cnt;

                if (input_axis_tlast) begin
                    status_valid_next = 1;
                    status_frame_pad_next = 0;
                    status_frame_truncate_next = 1;
                    status_frame_length_next = length_max;
                    status_frame_original_length_next = frame_ptr_next;
                    input_axis_tready_next = output_axis_tready_int_early & status_ready;
                    frame_ptr_next = 0;
                    state_next = STATE_IDLE;
                end else begin
                    state_next = STATE_TRUNCATE;
                end
            end else begin
                state_next = STATE_TRUNCATE;
            end
        end
    endcase
end

always @(posedge clk or posedge rst) begin
    if (rst) begin
        state_reg <= STATE_IDLE;
        frame_ptr_reg <= 0;
        input_axis_tready_reg <= 0;
        last_word_data_reg <= 0;
        last_word_keep_reg <= 0;
        last_cycle_tuser_reg <= 0;
        status_valid_reg <= 0;
        status_frame_pad_reg <= 0;
        status_frame_truncate_reg <= 0;
        status_frame_length_reg <= 0;
        status_frame_original_length_reg <= 0;
    end else begin
        state_reg <= state_next;

        frame_ptr_reg <= frame_ptr_next;

        input_axis_tready_reg <= input_axis_tready_next;

        last_cycle_tuser_reg <= last_cycle_tuser_next;

        status_valid_reg <= status_valid_next;
        status_frame_pad_reg <= status_frame_pad_next;
        status_frame_truncate_reg <= status_frame_truncate_next;
        status_frame_length_reg <= status_frame_length_next;
        status_frame_original_length_reg <= status_frame_original_length_next;

        if (store_last_word) begin
            last_word_data_reg <= output_axis_tdata_int;
            last_word_keep_reg <= output_axis_tkeep_int;
        end
    end
end

// output datapath logic
reg [DATA_WIDTH-1:0] output_axis_tdata_reg = 0;
reg [KEEP_WIDTH-1:0] output_axis_tkeep_reg = 0;
reg                  output_axis_tvalid_reg = 0;
reg                  output_axis_tlast_reg = 0;
reg                  output_axis_tuser_reg = 0;

reg [DATA_WIDTH-1:0] temp_axis_tdata_reg = 0;
reg [KEEP_WIDTH-1:0] temp_axis_tkeep_reg = 0;
reg                  temp_axis_tvalid_reg = 0;
reg                  temp_axis_tlast_reg = 0;
reg                  temp_axis_tuser_reg = 0;

assign output_axis_tdata = output_axis_tdata_reg;
assign output_axis_tkeep = output_axis_tkeep_reg;
assign output_axis_tvalid = output_axis_tvalid_reg;
assign output_axis_tlast = output_axis_tlast_reg;
assign output_axis_tuser = output_axis_tuser_reg;

// enable ready input next cycle if output is ready or if there is space in both output registers or if there is space in the temp register that will not be filled next cycle
assign output_axis_tready_int_early = output_axis_tready | (~temp_axis_tvalid_reg & ~output_axis_tvalid_reg) | (~temp_axis_tvalid_reg & ~output_axis_tvalid_int);

always @(posedge clk or posedge rst) begin
    if (rst) begin
        output_axis_tdata_reg <= 0;
        output_axis_tkeep_reg <= 0;
        output_axis_tvalid_reg <= 0;
        output_axis_tlast_reg <= 0;
        output_axis_tuser_reg <= 0;
        output_axis_tready_int <= 0;
        temp_axis_tdata_reg <= 0;
        temp_axis_tkeep_reg <= 0;
        temp_axis_tvalid_reg <= 0;
        temp_axis_tlast_reg <= 0;
        temp_axis_tuser_reg <= 0;
    end else begin
        // transfer sink ready state to source
        output_axis_tready_int <= output_axis_tready_int_early;

        if (output_axis_tready_int) begin
            // input is ready
            if (output_axis_tready | ~output_axis_tvalid_reg) begin
                // output is ready or currently not valid, transfer data to output
                output_axis_tdata_reg <= output_axis_tdata_int;
                output_axis_tkeep_reg <= output_axis_tkeep_int;
                output_axis_tvalid_reg <= output_axis_tvalid_int;
                output_axis_tlast_reg <= output_axis_tlast_int;
                output_axis_tuser_reg <= output_axis_tuser_int;
            end else begin
                // output is not ready and currently valid, store input in temp
                temp_axis_tdata_reg <= output_axis_tdata_int;
                temp_axis_tkeep_reg <= output_axis_tkeep_int;
                temp_axis_tvalid_reg <= output_axis_tvalid_int;
                temp_axis_tlast_reg <= output_axis_tlast_int;
                temp_axis_tuser_reg <= output_axis_tuser_int;
            end
        end else if (output_axis_tready) begin
            // input is not ready, but output is ready
            output_axis_tdata_reg <= temp_axis_tdata_reg;
            output_axis_tkeep_reg <= temp_axis_tkeep_reg;
            output_axis_tvalid_reg <= temp_axis_tvalid_reg;
            output_axis_tlast_reg <= temp_axis_tlast_reg;
            output_axis_tuser_reg <= temp_axis_tuser_reg;
            temp_axis_tdata_reg <= 0;
            temp_axis_tkeep_reg <= 0;
            temp_axis_tvalid_reg <= 0;
            temp_axis_tlast_reg <= 0;
            temp_axis_tuser_reg <= 0;
        end
    end
end

endmodule
