/*

Copyright (c) 2014-2016 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * Testbench for eth_demux_4
 */
module test_eth_demux_4;

// Inputs
reg clk = 0;
reg rst = 0;
reg [7:0] current_test = 0;

reg input_eth_hdr_valid = 0;
reg [47:0] input_eth_dest_mac = 0;
reg [47:0] input_eth_src_mac = 0;
reg [15:0] input_eth_type = 0;
reg [7:0] input_eth_payload_tdata = 0;
reg input_eth_payload_tvalid = 0;
reg input_eth_payload_tlast = 0;
reg input_eth_payload_tuser = 0;

reg output_0_eth_hdr_ready = 0;
reg output_0_eth_payload_tready = 0;
reg output_1_eth_hdr_ready = 0;
reg output_1_eth_payload_tready = 0;
reg output_2_eth_hdr_ready = 0;
reg output_2_eth_payload_tready = 0;
reg output_3_eth_hdr_ready = 0;
reg output_3_eth_payload_tready = 0;

reg enable = 0;
reg [1:0] select = 0;

// Outputs
wire input_eth_hdr_ready;
wire input_eth_payload_tready;

wire output_0_eth_hdr_valid;
wire [47:0] output_0_eth_dest_mac;
wire [47:0] output_0_eth_src_mac;
wire [15:0] output_0_eth_type;
wire [7:0] output_0_eth_payload_tdata;
wire output_0_eth_payload_tvalid;
wire output_0_eth_payload_tlast;
wire output_0_eth_payload_tuser;
wire output_1_eth_hdr_valid;
wire [47:0] output_1_eth_dest_mac;
wire [47:0] output_1_eth_src_mac;
wire [15:0] output_1_eth_type;
wire [7:0] output_1_eth_payload_tdata;
wire output_1_eth_payload_tvalid;
wire output_1_eth_payload_tlast;
wire output_1_eth_payload_tuser;
wire output_2_eth_hdr_valid;
wire [47:0] output_2_eth_dest_mac;
wire [47:0] output_2_eth_src_mac;
wire [15:0] output_2_eth_type;
wire [7:0] output_2_eth_payload_tdata;
wire output_2_eth_payload_tvalid;
wire output_2_eth_payload_tlast;
wire output_2_eth_payload_tuser;
wire output_3_eth_hdr_valid;
wire [47:0] output_3_eth_dest_mac;
wire [47:0] output_3_eth_src_mac;
wire [15:0] output_3_eth_type;
wire [7:0] output_3_eth_payload_tdata;
wire output_3_eth_payload_tvalid;
wire output_3_eth_payload_tlast;
wire output_3_eth_payload_tuser;

initial begin
    // myhdl integration
    $from_myhdl(
        clk,
        rst,
        current_test,
        input_eth_hdr_valid,
        input_eth_dest_mac,
        input_eth_src_mac,
        input_eth_type,
        input_eth_payload_tdata,
        input_eth_payload_tvalid,
        input_eth_payload_tlast,
        input_eth_payload_tuser,
        output_0_eth_hdr_ready,
        output_0_eth_payload_tready,
        output_1_eth_hdr_ready,
        output_1_eth_payload_tready,
        output_2_eth_hdr_ready,
        output_2_eth_payload_tready,
        output_3_eth_hdr_ready,
        output_3_eth_payload_tready,
        enable,
        select
    );
    $to_myhdl(
        input_eth_hdr_ready,
        input_eth_payload_tready,
        output_0_eth_hdr_valid,
        output_0_eth_dest_mac,
        output_0_eth_src_mac,
        output_0_eth_type,
        output_0_eth_payload_tdata,
        output_0_eth_payload_tvalid,
        output_0_eth_payload_tlast,
        output_0_eth_payload_tuser,
        output_1_eth_hdr_valid,
        output_1_eth_dest_mac,
        output_1_eth_src_mac,
        output_1_eth_type,
        output_1_eth_payload_tdata,
        output_1_eth_payload_tvalid,
        output_1_eth_payload_tlast,
        output_1_eth_payload_tuser,
        output_2_eth_hdr_valid,
        output_2_eth_dest_mac,
        output_2_eth_src_mac,
        output_2_eth_type,
        output_2_eth_payload_tdata,
        output_2_eth_payload_tvalid,
        output_2_eth_payload_tlast,
        output_2_eth_payload_tuser,
        output_3_eth_hdr_valid,
        output_3_eth_dest_mac,
        output_3_eth_src_mac,
        output_3_eth_type,
        output_3_eth_payload_tdata,
        output_3_eth_payload_tvalid,
        output_3_eth_payload_tlast,
        output_3_eth_payload_tuser
    );

    // dump file
    $dumpfile("test_eth_demux_4.lxt");
    $dumpvars(0, test_eth_demux_4);
end

eth_demux_4
UUT (
    .clk(clk),
    .rst(rst),
    // Ethernet frame input
    .input_eth_hdr_valid(input_eth_hdr_valid),
    .input_eth_hdr_ready(input_eth_hdr_ready),
    .input_eth_dest_mac(input_eth_dest_mac),
    .input_eth_src_mac(input_eth_src_mac),
    .input_eth_type(input_eth_type),
    .input_eth_payload_tdata(input_eth_payload_tdata),
    .input_eth_payload_tvalid(input_eth_payload_tvalid),
    .input_eth_payload_tready(input_eth_payload_tready),
    .input_eth_payload_tlast(input_eth_payload_tlast),
    .input_eth_payload_tuser(input_eth_payload_tuser),
    // Ethernet frame outputs
    .output_0_eth_hdr_valid(output_0_eth_hdr_valid),
    .output_0_eth_hdr_ready(output_0_eth_hdr_ready),
    .output_0_eth_dest_mac(output_0_eth_dest_mac),
    .output_0_eth_src_mac(output_0_eth_src_mac),
    .output_0_eth_type(output_0_eth_type),
    .output_0_eth_payload_tdata(output_0_eth_payload_tdata),
    .output_0_eth_payload_tvalid(output_0_eth_payload_tvalid),
    .output_0_eth_payload_tready(output_0_eth_payload_tready),
    .output_0_eth_payload_tlast(output_0_eth_payload_tlast),
    .output_0_eth_payload_tuser(output_0_eth_payload_tuser),
    .output_1_eth_hdr_valid(output_1_eth_hdr_valid),
    .output_1_eth_hdr_ready(output_1_eth_hdr_ready),
    .output_1_eth_dest_mac(output_1_eth_dest_mac),
    .output_1_eth_src_mac(output_1_eth_src_mac),
    .output_1_eth_type(output_1_eth_type),
    .output_1_eth_payload_tdata(output_1_eth_payload_tdata),
    .output_1_eth_payload_tvalid(output_1_eth_payload_tvalid),
    .output_1_eth_payload_tready(output_1_eth_payload_tready),
    .output_1_eth_payload_tlast(output_1_eth_payload_tlast),
    .output_1_eth_payload_tuser(output_1_eth_payload_tuser),
    .output_2_eth_hdr_valid(output_2_eth_hdr_valid),
    .output_2_eth_hdr_ready(output_2_eth_hdr_ready),
    .output_2_eth_dest_mac(output_2_eth_dest_mac),
    .output_2_eth_src_mac(output_2_eth_src_mac),
    .output_2_eth_type(output_2_eth_type),
    .output_2_eth_payload_tdata(output_2_eth_payload_tdata),
    .output_2_eth_payload_tvalid(output_2_eth_payload_tvalid),
    .output_2_eth_payload_tready(output_2_eth_payload_tready),
    .output_2_eth_payload_tlast(output_2_eth_payload_tlast),
    .output_2_eth_payload_tuser(output_2_eth_payload_tuser),
    .output_3_eth_hdr_valid(output_3_eth_hdr_valid),
    .output_3_eth_hdr_ready(output_3_eth_hdr_ready),
    .output_3_eth_dest_mac(output_3_eth_dest_mac),
    .output_3_eth_src_mac(output_3_eth_src_mac),
    .output_3_eth_type(output_3_eth_type),
    .output_3_eth_payload_tdata(output_3_eth_payload_tdata),
    .output_3_eth_payload_tvalid(output_3_eth_payload_tvalid),
    .output_3_eth_payload_tready(output_3_eth_payload_tready),
    .output_3_eth_payload_tlast(output_3_eth_payload_tlast),
    .output_3_eth_payload_tuser(output_3_eth_payload_tuser),
    // Control
    .enable(enable),
    .select(select)
);

endmodule
