/*

Copyright (c) 2014-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`timescale 1ns / 1ps

/*
 * LocalLink to AXI4-Stream bridge
 */
module ll_axis_bridge #
(
    parameter DATA_WIDTH = 8
)
(
    input  wire                   clk,
    input  wire                   rst,

    /*
     * LocalLink input
     */
    input  wire [DATA_WIDTH-1:0]  ll_data_in,
    input  wire                   ll_sof_in_n,
    input  wire                   ll_eof_in_n,
    input  wire                   ll_src_rdy_in_n,
    output wire                   ll_dst_rdy_out_n,

    /*
     * AXI output
     */
    output wire [DATA_WIDTH-1:0]  axis_tdata,
    output wire                   axis_tvalid,
    input  wire                   axis_tready,
    output wire                   axis_tlast
);

assign axis_tdata = ll_data_in;
assign axis_tvalid = ~ll_src_rdy_in_n;
assign axis_tlast = ~ll_eof_in_n;

assign ll_dst_rdy_out_n = ~axis_tready;

endmodule
